`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.09.2024 22:10:22
// Design Name: 
// Module Name: bit32_not
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:44:56 09/04/2024 
// Design Name: 
// Module Name:    bit8_not 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bit32_not(input wire [31:0] a,output wire [31:0] z);
not n0(z[0],a[0]);
not n1(z[1],a[1]);
not n2(z[2],a[2]);
not n3(z[3],a[3]);
not n4(z[4],a[4]);
not n5(z[5],a[5]);
not n6(z[6],a[6]);
not n7(z[7],a[7]);
not n8(z[8],a[8]);
not n9(z[9],a[9]);
not n10(z[10],a[10]);
not n11(z[11],a[11]);
not n12(z[12],a[12]);
not n13(z[13],a[13]);
not n14(z[14],a[14]);
not n15(z[15],a[15]);
not n16(z[16],a[16]);
not n17(z[17],a[17]);
not n18(z[18],a[18]);
not n19(z[19],a[19]);
not n20(z[20],a[20]);
not n21(z[21],a[21]);
not n22(z[22],a[22]);
not n23(z[23],a[23]);
not n24(z[24],a[24]);
not n25(z[25],a[25]);
not n26(z[26],a[26]);
not n27(z[27],a[27]);
not n28(z[28],a[28]);
not n29(z[29],a[29]);
not n30(z[30],a[30]);
not n31(z[31],a[31]);
endmodule
