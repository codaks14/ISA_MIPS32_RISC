`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04.11.2024 23:04:48
// Design Name: 
// Module Name: control_signal
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module control_signal(input wire optemp,input wire [5:0] func,input wire [4:0] opcode,input wire sloclock,output reg camehere,output reg load_PC,output reg load_IR,output reg select_MUX1,output reg select_MUX3,output reg select_MUX2,output reg select_MUX6,output reg write_REG,output reg [2:0] timesta,output reg select_MUX4,input rst,output reg [3:0] ALU_FUNC,output reg select_ALUOUT,output reg select_MUX5,output reg select_MUX7,output reg weaDM,output reg COMPout,output reg select_MUX8);

reg [2:0] next_state,state;


always @(state)
    case (state)
        3'b000:next_state<=3'b001;
        3'b001:next_state<=3'b010;
        3'b010:next_state<=3'b011;
        3'b011:next_state<=3'b100;
        3'b100:next_state<=3'b101;
        3'b101:next_state<=3'b110;
        default: next_state<=3'b000;
        endcase
        
always @(posedge sloclock)
    begin
    if(rst)
        begin
        load_IR=0;
        select_MUX1=0;
        select_MUX2=0;
        select_MUX3=0;
        select_MUX4=0;
        select_MUX6=0;
        write_REG=0;
        select_ALUOUT=0;
        timesta=0;
        load_PC=0;
        camehere=0;
        state<=3'b000;
        end
    else state<=next_state;
 end

localparam z4 = 4'b0000;
localparam ADD = 5'b00000;
localparam SUB = 5'b00001;
localparam AND = 5'b00010;
localparam OR = 5'b00011;
localparam XOR = 5'b00100;
localparam NOR = 5'b00101;
localparam NOT = 5'b00110;
localparam SL = 5'b00111;
localparam SRL = 5'b01000;
localparam SRA = 5'b01001;
localparam INC = 5'b01010;
localparam DEC = 5'b01011;
localparam SLT = 5'b01100;
localparam SGT = 5'b01101;
localparam HAM = 5'b01110;
localparam MOVE = 5'b01111;
localparam CMOV = 5'b10000;

localparam ADDI = 5'b00001;
localparam SUBI = 5'b00010;
localparam ANDI = 5'b00011;
localparam ORI = 5'b00100;
localparam XORI = 5'b00101;
localparam NORI = 5'b00110;
localparam NOTI = 5'b00111;
localparam SLAI = 5'b01000;
localparam SRLI = 5'b01001;
localparam SRAI = 5'b01010;
localparam SLTI = 5'b01011;
localparam SGTI = 5'b01100;
localparam HAMI = 5'b01101;
localparam LD = 5'b01110;
localparam ST = 5'b01111;
localparam BMI = 5'b10000;
localparam BPL = 5'b10001;
localparam BZ = 5'b10010;
localparam LUI = 5'b10011;
localparam BR = 5'b10100;
localparam HALT = 5'b10101;
localparam NOP = 5'b10110;

always @(state or opcode)
        begin
        if(opcode==5'b01111)begin
    if(state==0)
    begin
        load_PC<=0;
        load_IR<=1;
        write_REG<=0;
        select_MUX1<=0;
        select_MUX2<=0;
        select_MUX3<=0;
        select_MUX4<=0;
        select_MUX5<=0;
        select_MUX6<=0;
        select_MUX7<=0;
        select_MUX8<=0;
        select_ALUOUT<=0;
        ALU_FUNC<=4'b0000;
        weaDM<=0;  
    end
    else if(state==1)
    begin
        load_PC<=0;
        load_IR<=0;
        write_REG<=0;
        select_MUX1<=0;
        select_MUX2<=1;
        select_MUX3<=0;
        select_MUX4<=0;
        select_MUX5<=0;
        select_MUX6<=0;
        select_MUX7<=0;
        select_MUX8<=0;
        select_ALUOUT<=1;
        ALU_FUNC<=4'b0000;
        weaDM<=0;
    end
    else if(state==2)
    begin
        load_PC<=1;
        load_IR<=0;
        write_REG<=0;
        select_MUX1<=0;
        select_MUX2<=1;
        select_MUX3<=0;
        select_MUX4<=0;
        select_MUX5<=0;
        select_MUX6<=0;
        select_MUX7<=1;
        select_MUX8<=0;
        select_ALUOUT<=0;
        ALU_FUNC<=4'b0000;
        weaDM<=1; 
    end
//    if(state==3)
//    begin
//        load_PC<=1;
//        load_IR<=0;
//        write_REG<=0;
//        select_MUX1<=0;
//        select_MUX2<=0;
//        select_MUX3<=0;
//        select_MUX4<=0;
//        select_MUX5<=0;
//        select_MUX6<=0;
//        select_MUX7<=1;
//        select_MUX8<=0;
//        select_ALUOUT<=0;
//        ALU_FUNC<=4'b0000;
//        weaDM<=1;
//    end
    else 
    begin
        load_PC<=0;
        load_IR<=0;
        write_REG<=0;
        select_MUX1<=0;
        select_MUX2<=0;
        select_MUX3<=0;
        select_MUX4<=0;
        select_MUX5<=0;
        select_MUX6<=0;
        select_MUX7<=0;
        select_MUX8<=0;
        select_ALUOUT<=0;
        ALU_FUNC<=4'b0000;
        weaDM<=0;
    end
end
        if(optemp==0)
        begin
            if(func==ADD || func==SUB || func==AND || func==OR || func==XOR || func==NOR || func==NOT || func==SL || func==SRL || func==SRA || func==INC || func==DEC || func==SLT || func==SGT || func==HAM)
                begin
                    if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=1;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=func[3:0];
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                            select_MUX8<=0;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                     select_MUX8<=0;
                    end
                end
       end
       else
          begin
            if(opcode==ADDI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b0000;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end
            if(opcode==SUBI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=SUB;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end
            if(opcode==ANDI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b0010;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end

if(opcode==ORI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b0011;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end


if(opcode==XORI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b0100;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end

        
if(opcode==NORI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b0101;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end


if(opcode==NOTI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b0110;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end
          end
          if(opcode==SLAI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b0111;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end


if(opcode==SRLI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b1000;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end

if(opcode==SRAI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b1001;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end


if(opcode==SLTI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b1010;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end

if(opcode==SGTI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b1011;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end

if(opcode==HAMI)
            begin
                if(state==0)
                        begin
                            load_IR<=1;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            select_ALUOUT<=0;
                            select_MUX6<=0;
                            write_REG<=0;   
                            load_PC<=0;
                            select_MUX8<=0;
                            ALU_FUNC<=0;
                        end
                    else if(state==1)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_MUX2<=1;
                            select_MUX5<=0;
                            select_MUX7<=0;
                            ALU_FUNC<=4'b1100;
                            select_ALUOUT<=1;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=0;
                            load_PC<=0;
                            weaDM<=0; 
                            COMPout<=0;
                            select_MUX8<=0;
                        end
                    else if(state==2)
                        begin
                            load_IR<=0;
                            select_MUX1<=0;
                            select_MUX3<=0;
                            select_ALUOUT<=0;
                            select_MUX2<=0;
                            select_MUX4<=0;
                            select_MUX6<=0;
                            write_REG<=1;
                            load_PC<=1;
                            select_MUX5<=0;
                            select_MUX7<=1;
                            COMPout<=0;
                            weaDM<=0;
                            ALU_FUNC<=4'b0000;
                        end
                    else
                    begin
                     load_IR<=0;
                     select_MUX1<=0;
                     select_MUX3<=0;
                     select_MUX2<=0;
                     select_MUX4<=0;
                     select_MUX6<=0;
                     write_REG<=0;
                     load_PC<=0;
                     select_MUX5<=0;
                     select_MUX7<=0;
                     COMPout<=0;
                     weaDM<=0;
                     ALU_FUNC=4'b0000;
                    end
            end
if(opcode==BR)
    begin
        if(state==0)
            begin
                load_PC<=0;
                load_IR<=1;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=0;
                select_MUX8<=1;
                select_ALUOUT<=0;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
            else if(state==2)
            begin
                load_PC<=0;
                load_IR<=0;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=0;
                select_MUX8<=1;
                select_ALUOUT<=1;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
            else if(state==3)
            begin
                load_PC<=1;
                load_IR<=0;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=1;
                select_MUX8<=0;
                select_ALUOUT<=0;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
    end
if(opcode==BMI)
    begin
        if(state==0)
            begin
                load_PC<=0;
                load_IR<=1;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=0;
                select_MUX8<=0;
                select_ALUOUT<=0;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
            else if(state==2)
            begin
                load_PC<=0;
                load_IR<=0;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=0;
                select_MUX8<=0;
                select_ALUOUT<=1;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
            else if(state==3)
            begin
                load_PC<=1;
                load_IR<=0;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=1;
                select_MUX8<=0;
                select_ALUOUT<=0;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
    end
if(opcode==BPL)
    begin
        if(state==0)
            begin
                load_PC<=0;
                load_IR<=1;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=0;
                select_MUX8<=0;
                select_ALUOUT<=0;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
            else if(state==2)
            begin
                load_PC<=0;
                load_IR<=0;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=0;
                select_MUX8<=0;
                select_ALUOUT<=1;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
            else if(state==3)
            begin
                load_PC<=1;
                load_IR<=0;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=1;
                select_MUX8<=0;
                select_ALUOUT<=0;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
    end
if(opcode==BZ)
    begin
        if(state==0)
            begin
                load_PC<=0;
                load_IR<=1;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=0;
                select_MUX8<=0;
                select_ALUOUT<=0;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
            else if(state==2)
            begin
                load_PC<=0;
                load_IR<=0;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=0;
                select_MUX8<=0;
                select_ALUOUT<=1;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
            else if(state==3)
            begin
                load_PC<=1;
                load_IR<=0;
                write_REG<=0;
                select_MUX1<=0;
                select_MUX2<=0;
                select_MUX3<=0;
                select_MUX4<=0;
                select_MUX5<=0;
                select_MUX6<=0;
                select_MUX7<=1;
                select_MUX8<=0;
                select_ALUOUT<=0;
                ALU_FUNC<=4'b0000;
                weaDM<=0;
            end
    end
if(opcode==5'b01110)begin
    if(state==0)
    begin
        load_PC<=0;
        load_IR<=1;
        write_REG<=0;
        select_MUX1<=0;
        select_MUX2<=0;
        select_MUX3<=0;
        select_MUX4<=0;
        select_MUX5<=0;
        select_MUX6<=0;
        select_MUX7<=0;
        select_MUX8<=0;
        select_ALUOUT<=0;
        ALU_FUNC<=4'b0000;
        weaDM<=0;
       end   
       else if(state==1)
       begin
        load_PC<=0;
        load_IR<=0;
        write_REG<=0;
        select_MUX1<=0;
        select_MUX2<=1;
        select_MUX3<=0;
        select_MUX4<=0;
        select_MUX5<=0;
        select_MUX6<=0;
        select_MUX7<=0;
        select_MUX8<=0;
        select_ALUOUT<=1;
        ALU_FUNC<=4'b0000;
        weaDM<=0;
       end
       else if(state==2)
       begin
        load_PC<=1;
        load_IR<=0;
        write_REG<=1;
        select_MUX1<=0;
        select_MUX2<=0;
        select_MUX3<=0;
        select_MUX4<=0;
        select_MUX5<=0;
        select_MUX6<=0;
        select_MUX7<=1;
        select_MUX8<=0;
        select_ALUOUT<=0;
        ALU_FUNC<=4'b0000;
        weaDM<=0;
       end
       else
            begin
             load_IR<=0;
             select_MUX1<=0;
             select_MUX3<=0;
             select_MUX2<=0;
             select_MUX4<=0;
             select_MUX6<=0;
             write_REG<=0;
             load_PC<=0;
             select_MUX5<=0;
             select_MUX7<=0;
             COMPout<=0;
             weaDM<=0;
             ALU_FUNC=4'b0000;
            end
        end
if(opcode==5'b10101)
    begin
        if(state==1)
        begin
            load_PC<=0;
        end
    end
    end
endmodule
