`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.09.2024 18:50:46
// Design Name: 
// Module Name: bit32_leftshift
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bit32_leftshift(input wire [31:0] a,input wire [31:0] b,output wire [31:0] s);
wire [31:0] t;
mux32_1 b0(a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[0]);
mux32_1 b1(a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[1]);
mux32_1 b2(a[2],a[1],a[0],1'b0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[2]);
mux32_1 b3(a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[3]);
mux32_1 b4(a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[4]);
mux32_1 b5(a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[5]);
mux32_1 b6(a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[6]);
mux32_1 b7(a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[7]);
mux32_1 b8(a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[8]);
mux32_1 b9(a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[9]);
mux32_1 b10(a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[10]);
mux32_1 b11(a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[11]);
mux32_1 b12(a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[12]);
mux32_1 b13(a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[13]);
mux32_1 b14(a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[14]);
mux32_1 b15(a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[15]);
mux32_1 b16(a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[16]);
mux32_1 b17(a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[17]);
mux32_1 b18(a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[18]);
mux32_1 b19(a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[19]);
mux32_1 b20(a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,0,b[4:0],t[20]);
mux32_1 b21(a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,0,b[4:0],t[21]);
mux32_1 b22(a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,0,b[4:0],t[22]);
mux32_1 b23(a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,0,b[4:0],t[23]);
mux32_1 b24(a[24],a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,0,b[4:0],t[24]);
mux32_1 b25(a[25],a[24],a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,0,b[4:0],t[25]);
mux32_1 b26(a[26],a[25],a[24],a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,0,b[4:0],t[26]);
mux32_1 b27(a[27],a[26],a[25],a[24],a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,0,b[4:0],t[27]);
mux32_1 b28(a[28],a[27],a[26],a[25],a[24],a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,0,b[4:0],t[28]);
mux32_1 b29(a[29],a[28],a[27],a[26],a[25],a[24],a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,0,b[4:0],t[29]);
mux32_1 b30(a[30],a[29],a[28],a[27],a[26],a[25],a[24],a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],0,b[4:0],t[30]);
mux32_1 b31(a[31],a[30],a[29],a[28],a[27],a[26],a[25],a[24],a[23],a[22],a[21],a[20],a[19],a[18],a[17],a[16],a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0],b[4:0],t[31]);


or (e,b[5],b[6],b[7],b[8],b[9],b[10],b[11],b[12],b[13],b[14],b[15],b[16],b[17],b[18],b[19],b[20],b[21],b[22],b[23],b[24],b[25],b[26],b[27],b[28],b[29],b[30],b[31]);
Muxt2_1 m0(t,32'b0,e,s);
//assign s=t[31:0];


endmodule
